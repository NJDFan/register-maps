-- VHDL-2008 WISHBONE B4 package definitions.

package wishbone is
end package wishbone;

package body wishbone is
end package body wishbone;
